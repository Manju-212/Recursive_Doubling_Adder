//64 bit Recursive Doubling Adder
module Recursive_Doubling_Adder(A,B,Cin,Sum,Cout);

input [63:0] A,B;
output [64:0] Sum;input [1:0] Cin;
output Cout;

wire [1:0] kgp_0 [63:0];
wire [1:0] kgp_1 [63:0];
wire [1:0] kgp_2 [63:0];
wire [1:0] kgp_3 [63:0];
wire [1:0] kgp_4 [63:0];
wire [1:0] kgp_5 [63:0];
wire [1:0] kgp_6 [63:0];
wire [1:0] kgp_7 [63:0];
wire [1:0] kgp_8 [63:0];
wire [1:0] kgp_9 [63:0];
wire [1:0] kgp_10 [63:0];
wire [1:0] kgp_11 [63:0];
wire [1:0] kgp_12 [63:0];
wire [1:0] kgp_13 [63:0];
wire [1:0] kgp_14 [63:0];
wire [1:0] kgp_15 [63:0];
wire [1:0] kgp_16 [63:0];
wire [63:0] x_sum;


wire [64:0] carry;


assign carry[0] = Cin[0];

assign kgp_0[0]={A[0],B[0]};
assign kgp_0[1]={A[1],B[1]};
assign kgp_0[2]={A[2],B[2]};
assign kgp_0[3]={A[3],B[3]};
assign kgp_0[4]={A[4],B[4]};
assign kgp_0[5]={A[5],B[5]};
assign kgp_0[6]={A[6],B[6]};
assign kgp_0[7]={A[7],B[7]};
assign kgp_0[8]={A[8],B[8]};
assign kgp_0[9]={A[9],B[9]};
assign kgp_0[10]={A[10],B[10]};
assign kgp_0[11]={A[11],B[11]};
assign kgp_0[12]={A[12],B[12]};
assign kgp_0[13]={A[13],B[13]};
assign kgp_0[14]={A[14],B[14]};
assign kgp_0[15]={A[15],B[15]};
assign kgp_0[16]={A[16],B[16]};
assign kgp_0[17]={A[17],B[17]};
assign kgp_0[18]={A[18],B[18]};
assign kgp_0[19]={A[19],B[19]};
assign kgp_0[20]={A[20],B[20]};
assign kgp_0[21]={A[21],B[21]};
assign kgp_0[22]={A[22],B[22]};
assign kgp_0[23]={A[23],B[23]};
assign kgp_0[24]={A[24],B[24]};
assign kgp_0[25]={A[25],B[25]};
assign kgp_0[26]={A[26],B[26]};
assign kgp_0[27]={A[27],B[27]};
assign kgp_0[28]={A[28],B[28]};
assign kgp_0[29]={A[29],B[29]};
assign kgp_0[30]={A[30],B[30]};
assign kgp_0[31]={A[31],B[31]};
assign kgp_0[32]={A[32],B[32]};
assign kgp_0[33]={A[33],B[33]};
assign kgp_0[34]={A[34],B[34]};
assign kgp_0[35]={A[35],B[35]};
assign kgp_0[36]={A[36],B[36]};
assign kgp_0[37]={A[37],B[37]};
assign kgp_0[38]={A[38],B[38]};
assign kgp_0[39]={A[39],B[39]};
assign kgp_0[40]={A[40],B[40]};
assign kgp_0[41]={A[41],B[41]};
assign kgp_0[42]={A[42],B[42]};
assign kgp_0[43]={A[43],B[43]};
assign kgp_0[44]={A[44],B[44]};
assign kgp_0[45]={A[45],B[45]};
assign kgp_0[46]={A[46],B[46]};
assign kgp_0[47]={A[47],B[47]};
assign kgp_0[48]={A[48],B[48]};
assign kgp_0[49]={A[49],B[49]};
assign kgp_0[50]={A[50],B[50]};
assign kgp_0[51]={A[51],B[51]};
assign kgp_0[52]={A[52],B[52]};
assign kgp_0[53]={A[53],B[53]};
assign kgp_0[54]={A[54],B[54]};
assign kgp_0[55]={A[55],B[55]};
assign kgp_0[56]={A[56],B[56]};
assign kgp_0[57]={A[57],B[57]};
assign kgp_0[58]={A[58],B[58]};
assign kgp_0[59]={A[59],B[59]};
assign kgp_0[60]={A[60],B[60]};
assign kgp_0[61]={A[61],B[61]};
assign kgp_0[62]={A[62],B[62]};
assign kgp_0[63]={A[63],B[63]};



assign x_sum[0]=A[0]^B[0];
assign x_sum[1]=A[1]^B[1];
assign x_sum[2]=A[2]^B[2];
assign x_sum[3]=A[3]^B[3];
assign x_sum[4]=A[4]^B[4];
assign x_sum[5]=A[5]^B[5];
assign x_sum[6]=A[6]^B[6];
assign x_sum[7]=A[7]^B[7];
assign x_sum[8]=A[8]^B[8];
assign x_sum[9]=A[9]^B[9];
assign x_sum[10]=A[10]^B[10];
assign x_sum[11]=A[11]^B[11];
assign x_sum[12]=A[12]^B[12];
assign x_sum[13]=A[13]^B[13];
assign x_sum[14]=A[14]^B[14];
assign x_sum[15]=A[15]^B[15];
assign x_sum[16]=A[16]^B[16];
assign x_sum[17]=A[17]^B[17];
assign x_sum[18]=A[18]^B[18];
assign x_sum[19]=A[19]^B[19];
assign x_sum[20]=A[20]^B[20];
assign x_sum[21]=A[21]^B[21];
assign x_sum[22]=A[22]^B[22];
assign x_sum[23]=A[23]^B[23];
assign x_sum[24]=A[24]^B[24];
assign x_sum[25]=A[25]^B[25];
assign x_sum[26]=A[26]^B[26];
assign x_sum[27]=A[27]^B[27];
assign x_sum[28]=A[28]^B[28];
assign x_sum[29]=A[29]^B[29];
assign x_sum[30]=A[30]^B[30];
assign x_sum[31]=A[31]^B[31];
assign x_sum[32]=A[32]^B[32];
assign x_sum[33]=A[33]^B[33];
assign x_sum[34]=A[34]^B[34];
assign x_sum[35]=A[35]^B[35];
assign x_sum[36]=A[36]^B[36];
assign x_sum[37]=A[37]^B[37];
assign x_sum[38]=A[38]^B[38];
assign x_sum[39]=A[39]^B[39];
assign x_sum[40]=A[40]^B[40];
assign x_sum[41]=A[41]^B[41];
assign x_sum[42]=A[42]^B[42];
assign x_sum[43]=A[43]^B[43];
assign x_sum[44]=A[44]^B[44];
assign x_sum[45]=A[45]^B[45];
assign x_sum[46]=A[46]^B[46];
assign x_sum[47]=A[47]^B[47];
assign x_sum[48]=A[48]^B[48];
assign x_sum[49]=A[49]^B[49];
assign x_sum[50]=A[50]^B[50];
assign x_sum[51]=A[51]^B[51];
assign x_sum[52]=A[52]^B[52];
assign x_sum[53]=A[53]^B[53];
assign x_sum[54]=A[54]^B[54];
assign x_sum[55]=A[55]^B[55];
assign x_sum[56]=A[56]^B[56];
assign x_sum[57]=A[57]^B[57];
assign x_sum[58]=A[58]^B[58];
assign x_sum[59]=A[59]^B[59];
assign x_sum[60]=A[60]^B[60];
assign x_sum[61]=A[61]^B[61];
assign x_sum[62]=A[62]^B[62];
assign x_sum[63]=A[63]^B[63];

KGP k0(kgp_0[0],Cin,kgp_1[0]);
KGP k1(kgp_0[1],kgp_0[0],kgp_1[1]);
KGP k2(kgp_0[2],kgp_0[1],kgp_1[2]);
KGP k3(kgp_0[3],kgp_0[2],kgp_1[3]);
KGP k4(kgp_0[4],kgp_0[3],kgp_1[4]);
KGP k5(kgp_0[5],kgp_0[4],kgp_1[5]);
KGP k6(kgp_0[6],kgp_0[5],kgp_1[6]);
KGP k7(kgp_0[7],kgp_0[6],kgp_1[7]);
KGP k8(kgp_0[8],kgp_0[7],kgp_1[8]);
KGP k9(kgp_0[9],kgp_0[8],kgp_1[9]);
KGP k10(kgp_0[10],kgp_0[9],kgp_1[10]);
KGP k11(kgp_0[11],kgp_0[10],kgp_1[11]);
KGP k12(kgp_0[12],kgp_0[11],kgp_1[12]);
KGP k13(kgp_0[13],kgp_0[12],kgp_1[13]);
KGP k14(kgp_0[14],kgp_0[13],kgp_1[14]);
KGP k15(kgp_0[15],kgp_0[14],kgp_1[15]);
KGP k16(kgp_0[16],kgp_0[15],kgp_1[16]);
KGP k17(kgp_0[17],kgp_0[16],kgp_1[17]);
KGP k18(kgp_0[18],kgp_0[17],kgp_1[18]);
KGP k19(kgp_0[19],kgp_0[18],kgp_1[19]);
KGP k20(kgp_0[20],kgp_0[19],kgp_1[20]);
KGP k21(kgp_0[21],kgp_0[20],kgp_1[21]);
KGP k22(kgp_0[22],kgp_0[21],kgp_1[22]);
KGP k23(kgp_0[23],kgp_0[22],kgp_1[23]);
KGP k24(kgp_0[24],kgp_0[23],kgp_1[24]);
KGP k25(kgp_0[25],kgp_0[24],kgp_1[25]);
KGP k26(kgp_0[26],kgp_0[25],kgp_1[26]);
KGP k27(kgp_0[27],kgp_0[26],kgp_1[27]);
KGP k28(kgp_0[28],kgp_0[27],kgp_1[28]);
KGP k29(kgp_0[29],kgp_0[28],kgp_1[29]);
KGP k30(kgp_0[30],kgp_0[29],kgp_1[30]);
KGP k31(kgp_0[31],kgp_0[30],kgp_1[31]);
KGP k32(kgp_0[32],kgp_0[31],kgp_1[32]);
KGP k33(kgp_0[33],kgp_0[32],kgp_1[33]);
KGP k34(kgp_0[34],kgp_0[33],kgp_1[34]);
KGP k35(kgp_0[35],kgp_0[34],kgp_1[35]);
KGP k36(kgp_0[36],kgp_0[35],kgp_1[36]);
KGP k37(kgp_0[37],kgp_0[36],kgp_1[37]);
KGP k38(kgp_0[38],kgp_0[37],kgp_1[38]);
KGP k39(kgp_0[39],kgp_0[38],kgp_1[39]);
KGP k40(kgp_0[40],kgp_0[39],kgp_1[40]);
KGP k41(kgp_0[41],kgp_0[40],kgp_1[41]);
KGP k42(kgp_0[42],kgp_0[41],kgp_1[42]);
KGP k43(kgp_0[43],kgp_0[42],kgp_1[43]);
KGP k44(kgp_0[44],kgp_0[43],kgp_1[44]);
KGP k45(kgp_0[45],kgp_0[44],kgp_1[45]);
KGP k46(kgp_0[46],kgp_0[45],kgp_1[46]);
KGP k47(kgp_0[47],kgp_0[46],kgp_1[47]);
KGP k48(kgp_0[48],kgp_0[47],kgp_1[48]);
KGP k49(kgp_0[49],kgp_0[48],kgp_1[49]);
KGP k50(kgp_0[50],kgp_0[49],kgp_1[50]);
KGP k51(kgp_0[51],kgp_0[50],kgp_1[51]);
KGP k52(kgp_0[52],kgp_0[51],kgp_1[52]);
KGP k53(kgp_0[53],kgp_0[52],kgp_1[53]);
KGP k54(kgp_0[54],kgp_0[53],kgp_1[54]);
KGP k55(kgp_0[55],kgp_0[54],kgp_1[55]);
KGP k56(kgp_0[56],kgp_0[55],kgp_1[56]);
KGP k57(kgp_0[57],kgp_0[56],kgp_1[57]);
KGP k58(kgp_0[58],kgp_0[57],kgp_1[58]);
KGP k59(kgp_0[59],kgp_0[58],kgp_1[59]);
KGP k60(kgp_0[60],kgp_0[59],kgp_1[60]);
KGP k61(kgp_0[61],kgp_0[60],kgp_1[61]);
KGP k62(kgp_0[62],kgp_0[61],kgp_1[62]);
KGP k63(kgp_0[63],kgp_0[62],kgp_1[63]);



KGP k64(kgp_1[1],Cin,kgp_2[1]);
KGP k65(kgp_1[2],kgp_1[0],kgp_2[2]);
KGP k66(kgp_1[3],kgp_1[1],kgp_2[3]);
KGP k67(kgp_1[4],kgp_1[2],kgp_2[4]);
KGP k68(kgp_1[5],kgp_1[3],kgp_2[5]);
KGP k69(kgp_1[6],kgp_1[4],kgp_2[6]);
KGP k70(kgp_1[7],kgp_1[5],kgp_2[7]);
KGP k71(kgp_1[8],kgp_1[6],kgp_2[8]);
KGP k72(kgp_1[9],kgp_1[7],kgp_2[9]);
KGP k73(kgp_1[10],kgp_1[8],kgp_2[10]);
KGP k74(kgp_1[11],kgp_1[9],kgp_2[11]);
KGP k75(kgp_1[12],kgp_1[10],kgp_2[12]);
KGP k76(kgp_1[13],kgp_1[11],kgp_2[13]);
KGP k77(kgp_1[14],kgp_1[12],kgp_2[14]);
KGP k78(kgp_1[15],kgp_1[13],kgp_2[15]);
KGP k79(kgp_1[16],kgp_1[14],kgp_2[16]);
KGP k80(kgp_1[17],kgp_1[15],kgp_2[17]);
KGP k81(kgp_1[18],kgp_1[16],kgp_2[18]);
KGP k82(kgp_1[19],kgp_1[17],kgp_2[19]);
KGP k83(kgp_1[20],kgp_1[18],kgp_2[20]);
KGP k84(kgp_1[21],kgp_1[19],kgp_2[21]);
KGP k85(kgp_1[22],kgp_1[20],kgp_2[22]);
KGP k86(kgp_1[23],kgp_1[21],kgp_2[23]);
KGP k87(kgp_1[24],kgp_1[22],kgp_2[24]);
KGP k88(kgp_1[25],kgp_1[23],kgp_2[25]);
KGP k89(kgp_1[26],kgp_1[24],kgp_2[26]);
KGP k90(kgp_1[27],kgp_1[25],kgp_2[27]);
KGP k91(kgp_1[28],kgp_1[26],kgp_2[28]);
KGP k92(kgp_1[29],kgp_1[27],kgp_2[29]);
KGP k93(kgp_1[30],kgp_1[28],kgp_2[30]);
KGP k94(kgp_1[31],kgp_1[29],kgp_2[31]);
KGP k95(kgp_1[32],kgp_1[30],kgp_2[32]);
KGP k96(kgp_1[33],kgp_1[31],kgp_2[33]);
KGP k97(kgp_1[34],kgp_1[32],kgp_2[34]);
KGP k98(kgp_1[35],kgp_1[33],kgp_2[35]);
KGP k99(kgp_1[36],kgp_1[34],kgp_2[36]);
KGP k100(kgp_1[37],kgp_1[35],kgp_2[37]);
KGP k101(kgp_1[38],kgp_1[36],kgp_2[38]);
KGP k102(kgp_1[39],kgp_1[37],kgp_2[39]);
KGP k103(kgp_1[40],kgp_1[38],kgp_2[40]);
KGP k104(kgp_1[41],kgp_1[39],kgp_2[41]);
KGP k105(kgp_1[42],kgp_1[40],kgp_2[42]);
KGP k106(kgp_1[43],kgp_1[41],kgp_2[43]);
KGP k107(kgp_1[44],kgp_1[42],kgp_2[44]);
KGP k108(kgp_1[45],kgp_1[43],kgp_2[45]);
KGP k109(kgp_1[46],kgp_1[44],kgp_2[46]);
KGP k110(kgp_1[47],kgp_1[45],kgp_2[47]);
KGP k111(kgp_1[48],kgp_1[46],kgp_2[48]);
KGP k112(kgp_1[49],kgp_1[47],kgp_2[49]);
KGP k113(kgp_1[50],kgp_1[48],kgp_2[50]);
KGP k114(kgp_1[51],kgp_1[49],kgp_2[51]);
KGP k115(kgp_1[52],kgp_1[50],kgp_2[52]);
KGP k116(kgp_1[53],kgp_1[51],kgp_2[53]);
KGP k117(kgp_1[54],kgp_1[52],kgp_2[54]);
KGP k118(kgp_1[55],kgp_1[53],kgp_2[55]);
KGP k119(kgp_1[56],kgp_1[54],kgp_2[56]);
KGP k120(kgp_1[57],kgp_1[55],kgp_2[57]);
KGP k121(kgp_1[58],kgp_1[56],kgp_2[58]);
KGP k122(kgp_1[59],kgp_1[57],kgp_2[59]);
KGP k123(kgp_1[60],kgp_1[58],kgp_2[60]);
KGP k124(kgp_1[61],kgp_1[59],kgp_2[61]);
KGP k125(kgp_1[62],kgp_1[60],kgp_2[62]);
KGP k126(kgp_1[63],kgp_1[61],kgp_2[63]);



KGP k127(kgp_2[3],Cin,kgp_3[3]);
KGP k128(kgp_2[4],kgp_2[0],kgp_3[4]);
KGP k129(kgp_2[5],kgp_2[1],kgp_3[5]);
KGP k130(kgp_2[6],kgp_2[2],kgp_3[6]);
KGP k131(kgp_2[7],kgp_2[3],kgp_3[7]);
KGP k132(kgp_2[8],kgp_2[4],kgp_3[8]);
KGP k133(kgp_2[9],kgp_2[5],kgp_3[9]);
KGP k134(kgp_2[10],kgp_2[6],kgp_3[10]);
KGP k135(kgp_2[11],kgp_2[7],kgp_3[11]);
KGP k136(kgp_2[12],kgp_2[8],kgp_3[12]);
KGP k137(kgp_2[13],kgp_2[9],kgp_3[13]);
KGP k138(kgp_2[14],kgp_2[10],kgp_3[14]);
KGP k139(kgp_2[15],kgp_2[11],kgp_3[15]);
KGP k140(kgp_2[16],kgp_2[12],kgp_3[16]);
KGP k141(kgp_2[17],kgp_2[13],kgp_3[17]);
KGP k142(kgp_2[18],kgp_2[14],kgp_3[18]);
KGP k143(kgp_2[19],kgp_2[15],kgp_3[19]);
KGP k144(kgp_2[20],kgp_2[16],kgp_3[20]);
KGP k145(kgp_2[21],kgp_2[17],kgp_3[21]);
KGP k146(kgp_2[22],kgp_2[18],kgp_3[22]);
KGP k147(kgp_2[23],kgp_2[19],kgp_3[23]);
KGP k148(kgp_2[24],kgp_2[20],kgp_3[24]);
KGP k149(kgp_2[25],kgp_2[21],kgp_3[25]);
KGP k150(kgp_2[26],kgp_2[22],kgp_3[26]);
KGP k151(kgp_2[27],kgp_2[23],kgp_3[27]);
KGP k152(kgp_2[28],kgp_2[24],kgp_3[28]);
KGP k153(kgp_2[29],kgp_2[25],kgp_3[29]);
KGP k154(kgp_2[30],kgp_2[26],kgp_3[30]);
KGP k155(kgp_2[31],kgp_2[27],kgp_3[31]);
KGP k156(kgp_2[32],kgp_2[28],kgp_3[32]);
KGP k157(kgp_2[33],kgp_2[29],kgp_3[33]);
KGP k158(kgp_2[34],kgp_2[30],kgp_3[34]);
KGP k159(kgp_2[35],kgp_2[31],kgp_3[35]);
KGP k160(kgp_2[36],kgp_2[32],kgp_3[36]);
KGP k161(kgp_2[37],kgp_2[33],kgp_3[37]);
KGP k162(kgp_2[38],kgp_2[34],kgp_3[38]);
KGP k163(kgp_2[39],kgp_2[35],kgp_3[39]);
KGP k164(kgp_2[40],kgp_2[36],kgp_3[40]);
KGP k165(kgp_2[41],kgp_2[37],kgp_3[41]);
KGP k166(kgp_2[42],kgp_2[38],kgp_3[42]);
KGP k167(kgp_2[43],kgp_2[39],kgp_3[43]);
KGP k168(kgp_2[44],kgp_2[40],kgp_3[44]);
KGP k169(kgp_2[45],kgp_2[41],kgp_3[45]);
KGP k170(kgp_2[46],kgp_2[42],kgp_3[46]);
KGP k171(kgp_2[47],kgp_2[43],kgp_3[47]);
KGP k172(kgp_2[48],kgp_2[44],kgp_3[48]);
KGP k173(kgp_2[49],kgp_2[45],kgp_3[49]);
KGP k174(kgp_2[50],kgp_2[46],kgp_3[50]);
KGP k175(kgp_2[51],kgp_2[47],kgp_3[51]);
KGP k176(kgp_2[52],kgp_2[48],kgp_3[52]);
KGP k177(kgp_2[53],kgp_2[49],kgp_3[53]);
KGP k178(kgp_2[54],kgp_2[50],kgp_3[54]);
KGP k179(kgp_2[55],kgp_2[51],kgp_3[55]);
KGP k180(kgp_2[56],kgp_2[52],kgp_3[56]);
KGP k181(kgp_2[57],kgp_2[53],kgp_3[57]);
KGP k182(kgp_2[58],kgp_2[54],kgp_3[58]);
KGP k183(kgp_2[59],kgp_2[55],kgp_3[59]);
KGP k184(kgp_2[60],kgp_2[56],kgp_3[60]);
KGP k185(kgp_2[61],kgp_2[57],kgp_3[61]);
KGP k186(kgp_2[62],kgp_2[58],kgp_3[62]);
KGP k187(kgp_2[63],kgp_2[59],kgp_3[63]);



KGP k188(kgp_3[7],Cin,kgp_4[7]);
KGP k189(kgp_3[8],kgp_3[0],kgp_4[8]);
KGP k190(kgp_3[9],kgp_3[1],kgp_4[9]);
KGP k191(kgp_3[10],kgp_3[2],kgp_4[10]);
KGP k192(kgp_3[11],kgp_3[3],kgp_4[11]);
KGP k193(kgp_3[12],kgp_3[4],kgp_4[12]);
KGP k194(kgp_3[13],kgp_3[5],kgp_4[13]);
KGP k195(kgp_3[14],kgp_3[6],kgp_4[14]);
KGP k196(kgp_3[15],kgp_3[7],kgp_4[15]);
KGP k197(kgp_3[16],kgp_3[8],kgp_4[16]);
KGP k198(kgp_3[17],kgp_3[9],kgp_4[17]);
KGP k199(kgp_3[18],kgp_3[10],kgp_4[18]);
KGP k200(kgp_3[19],kgp_3[11],kgp_4[19]);
KGP k201(kgp_3[20],kgp_3[12],kgp_4[20]);
KGP k202(kgp_3[21],kgp_3[13],kgp_4[21]);
KGP k203(kgp_3[22],kgp_3[14],kgp_4[22]);
KGP k204(kgp_3[23],kgp_3[15],kgp_4[23]);
KGP k205(kgp_3[24],kgp_3[16],kgp_4[24]);
KGP k206(kgp_3[25],kgp_3[17],kgp_4[25]);
KGP k207(kgp_3[26],kgp_3[18],kgp_4[26]);
KGP k208(kgp_3[27],kgp_3[19],kgp_4[27]);
KGP k209(kgp_3[28],kgp_3[20],kgp_4[28]);
KGP k210(kgp_3[29],kgp_3[21],kgp_4[29]);
KGP k211(kgp_3[30],kgp_3[22],kgp_4[30]);
KGP k212(kgp_3[31],kgp_3[23],kgp_4[31]);
KGP k213(kgp_3[32],kgp_3[24],kgp_4[32]);
KGP k214(kgp_3[33],kgp_3[25],kgp_4[33]);
KGP k215(kgp_3[34],kgp_3[26],kgp_4[34]);
KGP k216(kgp_3[35],kgp_3[27],kgp_4[35]);
KGP k217(kgp_3[36],kgp_3[28],kgp_4[36]);
KGP k218(kgp_3[37],kgp_3[29],kgp_4[37]);
KGP k219(kgp_3[38],kgp_3[30],kgp_4[38]);
KGP k220(kgp_3[39],kgp_3[31],kgp_4[39]);
KGP k221(kgp_3[40],kgp_3[32],kgp_4[40]);
KGP k222(kgp_3[41],kgp_3[33],kgp_4[41]);
KGP k223(kgp_3[42],kgp_3[34],kgp_4[42]);
KGP k224(kgp_3[43],kgp_3[35],kgp_4[43]);
KGP k225(kgp_3[44],kgp_3[36],kgp_4[44]);
KGP k226(kgp_3[45],kgp_3[37],kgp_4[45]);
KGP k227(kgp_3[46],kgp_3[38],kgp_4[46]);
KGP k228(kgp_3[47],kgp_3[39],kgp_4[47]);
KGP k229(kgp_3[48],kgp_3[40],kgp_4[48]);
KGP k230(kgp_3[49],kgp_3[41],kgp_4[49]);
KGP k231(kgp_3[50],kgp_3[42],kgp_4[50]);
KGP k232(kgp_3[51],kgp_3[43],kgp_4[51]);
KGP k233(kgp_3[52],kgp_3[44],kgp_4[52]);
KGP k234(kgp_3[53],kgp_3[45],kgp_4[53]);
KGP k235(kgp_3[54],kgp_3[46],kgp_4[54]);
KGP k236(kgp_3[55],kgp_3[47],kgp_4[55]);
KGP k237(kgp_3[56],kgp_3[48],kgp_4[56]);
KGP k238(kgp_3[57],kgp_3[49],kgp_4[57]);
KGP k239(kgp_3[58],kgp_3[50],kgp_4[58]);
KGP k240(kgp_3[59],kgp_3[51],kgp_4[59]);
KGP k241(kgp_3[60],kgp_3[52],kgp_4[60]);
KGP k242(kgp_3[61],kgp_3[53],kgp_4[61]);
KGP k243(kgp_3[62],kgp_3[54],kgp_4[62]);
KGP k244(kgp_3[63],kgp_3[55],kgp_4[63]);



KGP k245(kgp_4[15],Cin,kgp_5[15]);
KGP k246(kgp_4[16],kgp_4[0],kgp_5[16]);
KGP k247(kgp_4[17],kgp_4[1],kgp_5[17]);
KGP k248(kgp_4[18],kgp_4[2],kgp_5[18]);
KGP k249(kgp_4[19],kgp_4[3],kgp_5[19]);
KGP k250(kgp_4[20],kgp_4[4],kgp_5[20]);
KGP k251(kgp_4[21],kgp_4[5],kgp_5[21]);
KGP k252(kgp_4[22],kgp_4[6],kgp_5[22]);
KGP k253(kgp_4[23],kgp_4[7],kgp_5[23]);
KGP k254(kgp_4[24],kgp_4[8],kgp_5[24]);
KGP k255(kgp_4[25],kgp_4[9],kgp_5[25]);
KGP k256(kgp_4[26],kgp_4[10],kgp_5[26]);
KGP k257(kgp_4[27],kgp_4[11],kgp_5[27]);
KGP k258(kgp_4[28],kgp_4[12],kgp_5[28]);
KGP k259(kgp_4[29],kgp_4[13],kgp_5[29]);
KGP k260(kgp_4[30],kgp_4[14],kgp_5[30]);
KGP k261(kgp_4[31],kgp_4[15],kgp_5[31]);
KGP k262(kgp_4[32],kgp_4[16],kgp_5[32]);
KGP k263(kgp_4[33],kgp_4[17],kgp_5[33]);
KGP k264(kgp_4[34],kgp_4[18],kgp_5[34]);
KGP k265(kgp_4[35],kgp_4[19],kgp_5[35]);
KGP k266(kgp_4[36],kgp_4[20],kgp_5[36]);
KGP k267(kgp_4[37],kgp_4[21],kgp_5[37]);
KGP k268(kgp_4[38],kgp_4[22],kgp_5[38]);
KGP k269(kgp_4[39],kgp_4[23],kgp_5[39]);
KGP k270(kgp_4[40],kgp_4[24],kgp_5[40]);
KGP k271(kgp_4[41],kgp_4[25],kgp_5[41]);
KGP k272(kgp_4[42],kgp_4[26],kgp_5[42]);
KGP k273(kgp_4[43],kgp_4[27],kgp_5[43]);
KGP k274(kgp_4[44],kgp_4[28],kgp_5[44]);
KGP k275(kgp_4[45],kgp_4[29],kgp_5[45]);
KGP k276(kgp_4[46],kgp_4[30],kgp_5[46]);
KGP k277(kgp_4[47],kgp_4[31],kgp_5[47]);
KGP k278(kgp_4[48],kgp_4[32],kgp_5[48]);
KGP k279(kgp_4[49],kgp_4[33],kgp_5[49]);
KGP k280(kgp_4[50],kgp_4[34],kgp_5[50]);
KGP k281(kgp_4[51],kgp_4[35],kgp_5[51]);
KGP k282(kgp_4[52],kgp_4[36],kgp_5[52]);
KGP k283(kgp_4[53],kgp_4[37],kgp_5[53]);
KGP k284(kgp_4[54],kgp_4[38],kgp_5[54]);
KGP k285(kgp_4[55],kgp_4[39],kgp_5[55]);
KGP k286(kgp_4[56],kgp_4[40],kgp_5[56]);
KGP k287(kgp_4[57],kgp_4[41],kgp_5[57]);
KGP k288(kgp_4[58],kgp_4[42],kgp_5[58]);
KGP k289(kgp_4[59],kgp_4[43],kgp_5[59]);
KGP k290(kgp_4[60],kgp_4[44],kgp_5[60]);
KGP k291(kgp_4[61],kgp_4[45],kgp_5[61]);
KGP k292(kgp_4[62],kgp_4[46],kgp_5[62]);
KGP k293(kgp_4[63],kgp_4[47],kgp_5[63]);



KGP k294(kgp_5[31],Cin,kgp_6[31]);
KGP k295(kgp_5[32],kgp_5[0],kgp_6[32]);
KGP k296(kgp_5[33],kgp_5[1],kgp_6[33]);
KGP k297(kgp_5[34],kgp_5[2],kgp_6[34]);
KGP k298(kgp_5[35],kgp_5[3],kgp_6[35]);
KGP k299(kgp_5[36],kgp_5[4],kgp_6[36]);
KGP k300(kgp_5[37],kgp_5[5],kgp_6[37]);
KGP k301(kgp_5[38],kgp_5[6],kgp_6[38]);
KGP k302(kgp_5[39],kgp_5[7],kgp_6[39]);
KGP k303(kgp_5[40],kgp_5[8],kgp_6[40]);
KGP k304(kgp_5[41],kgp_5[9],kgp_6[41]);
KGP k305(kgp_5[42],kgp_5[10],kgp_6[42]);
KGP k306(kgp_5[43],kgp_5[11],kgp_6[43]);
KGP k307(kgp_5[44],kgp_5[12],kgp_6[44]);
KGP k308(kgp_5[45],kgp_5[13],kgp_6[45]);
KGP k309(kgp_5[46],kgp_5[14],kgp_6[46]);
KGP k310(kgp_5[47],kgp_5[15],kgp_6[47]);
KGP k311(kgp_5[48],kgp_5[16],kgp_6[48]);
KGP k312(kgp_5[49],kgp_5[17],kgp_6[49]);
KGP k313(kgp_5[50],kgp_5[18],kgp_6[50]);
KGP k314(kgp_5[51],kgp_5[19],kgp_6[51]);
KGP k315(kgp_5[52],kgp_5[20],kgp_6[52]);
KGP k316(kgp_5[53],kgp_5[21],kgp_6[53]);
KGP k317(kgp_5[54],kgp_5[22],kgp_6[54]);
KGP k318(kgp_5[55],kgp_5[23],kgp_6[55]);
KGP k319(kgp_5[56],kgp_5[24],kgp_6[56]);
KGP k320(kgp_5[57],kgp_5[25],kgp_6[57]);
KGP k321(kgp_5[58],kgp_5[26],kgp_6[58]);
KGP k322(kgp_5[59],kgp_5[27],kgp_6[59]);
KGP k323(kgp_5[60],kgp_5[28],kgp_6[60]);
KGP k324(kgp_5[61],kgp_5[29],kgp_6[61]);
KGP k325(kgp_5[62],kgp_5[30],kgp_6[62]);
KGP k326(kgp_5[63],kgp_5[31],kgp_6[63]);



KGP k327(kgp_6[63],Cin,kgp_7[63]);




assign carry[1] = kgp_1[0][0];
assign carry[2] = kgp_2[1][0];
assign carry[3] = kgp_2[2][0];
assign carry[4] = kgp_2[3][0];
assign carry[5] = kgp_3[4][0];
assign carry[6] = kgp_3[5][0];
assign carry[7] = kgp_3[6][0];
assign carry[8] = kgp_3[7][0];
assign carry[9] = kgp_3[8][0];
assign carry[10] = kgp_3[9][0];
assign carry[11] = kgp_3[10][0];
assign carry[12] = kgp_4[11][0];
assign carry[13] = kgp_4[12][0];
assign carry[14] = kgp_4[13][0];
assign carry[15] = kgp_4[14][0];
assign carry[16] = kgp_4[15][0];
assign carry[17] = kgp_4[16][0];
assign carry[18] = kgp_4[17][0];
assign carry[19] = kgp_4[18][0];
assign carry[20] = kgp_4[19][0];
assign carry[21] = kgp_4[20][0];
assign carry[22] = kgp_4[21][0];
assign carry[23] = kgp_4[22][0];
assign carry[24] = kgp_4[23][0];
assign carry[25] = kgp_4[24][0];
assign carry[26] = kgp_4[25][0];
assign carry[27] = kgp_5[26][0];
assign carry[28] = kgp_5[27][0];
assign carry[29] = kgp_5[28][0];
assign carry[30] = kgp_5[29][0];
assign carry[31] = kgp_5[30][0];
assign carry[32] = kgp_5[31][0];
assign carry[33] = kgp_5[32][0];
assign carry[34] = kgp_5[33][0];
assign carry[35] = kgp_5[34][0];
assign carry[36] = kgp_5[35][0];
assign carry[37] = kgp_5[36][0];
assign carry[38] = kgp_5[37][0];
assign carry[39] = kgp_5[38][0];
assign carry[40] = kgp_5[39][0];
assign carry[41] = kgp_5[40][0];
assign carry[42] = kgp_5[41][0];
assign carry[43] = kgp_5[42][0];
assign carry[44] = kgp_5[43][0];
assign carry[45] = kgp_5[44][0];
assign carry[46] = kgp_5[45][0];
assign carry[47] = kgp_5[46][0];
assign carry[48] = kgp_5[47][0];
assign carry[49] = kgp_5[48][0];
assign carry[50] = kgp_5[49][0];
assign carry[51] = kgp_5[50][0];
assign carry[52] = kgp_5[51][0];
assign carry[53] = kgp_5[52][0];
assign carry[54] = kgp_5[53][0];
assign carry[55] = kgp_5[54][0];
assign carry[56] = kgp_5[55][0];
assign carry[57] = kgp_5[56][0];
assign carry[58] = kgp_6[57][0];
assign carry[59] = kgp_6[58][0];
assign carry[60] = kgp_6[59][0];
assign carry[61] = kgp_6[60][0];
assign carry[62] = kgp_6[61][0];
assign carry[63] = kgp_6[62][0];
assign carry[64] = kgp_6[63][0];
assign Cout = carry[64];

assign Sum[0]= x_sum[0] ^carry[0];
assign Sum[1]= x_sum[1] ^carry[1];
assign Sum[2]= x_sum[2] ^carry[2];
assign Sum[3]= x_sum[3] ^carry[3];
assign Sum[4]= x_sum[4] ^carry[4];
assign Sum[5]= x_sum[5] ^carry[5];
assign Sum[6]= x_sum[6] ^carry[6];
assign Sum[7]= x_sum[7] ^carry[7];
assign Sum[8]= x_sum[8] ^carry[8];
assign Sum[9]= x_sum[9] ^carry[9];
assign Sum[10]= x_sum[10] ^carry[10];
assign Sum[11]= x_sum[11] ^carry[11];
assign Sum[12]= x_sum[12] ^carry[12];
assign Sum[13]= x_sum[13] ^carry[13];
assign Sum[14]= x_sum[14] ^carry[14];
assign Sum[15]= x_sum[15] ^carry[15];
assign Sum[16]= x_sum[16] ^carry[16];
assign Sum[17]= x_sum[17] ^carry[17];
assign Sum[18]= x_sum[18] ^carry[18];
assign Sum[19]= x_sum[19] ^carry[19];
assign Sum[20]= x_sum[20] ^carry[20];
assign Sum[21]= x_sum[21] ^carry[21];
assign Sum[22]= x_sum[22] ^carry[22];
assign Sum[23]= x_sum[23] ^carry[23];
assign Sum[24]= x_sum[24] ^carry[24];
assign Sum[25]= x_sum[25] ^carry[25];
assign Sum[26]= x_sum[26] ^carry[26];
assign Sum[27]= x_sum[27] ^carry[27];
assign Sum[28]= x_sum[28] ^carry[28];
assign Sum[29]= x_sum[29] ^carry[29];
assign Sum[30]= x_sum[30] ^carry[30];
assign Sum[31]= x_sum[31] ^carry[31];
assign Sum[32]= x_sum[32] ^carry[32];
assign Sum[33]= x_sum[33] ^carry[33];
assign Sum[34]= x_sum[34] ^carry[34];
assign Sum[35]= x_sum[35] ^carry[35];
assign Sum[36]= x_sum[36] ^carry[36];
assign Sum[37]= x_sum[37] ^carry[37];
assign Sum[38]= x_sum[38] ^carry[38];
assign Sum[39]= x_sum[39] ^carry[39];
assign Sum[40]= x_sum[40] ^carry[40];
assign Sum[41]= x_sum[41] ^carry[41];
assign Sum[42]= x_sum[42] ^carry[42];
assign Sum[43]= x_sum[43] ^carry[43];
assign Sum[44]= x_sum[44] ^carry[44];
assign Sum[45]= x_sum[45] ^carry[45];
assign Sum[46]= x_sum[46] ^carry[46];
assign Sum[47]= x_sum[47] ^carry[47];
assign Sum[48]= x_sum[48] ^carry[48];
assign Sum[49]= x_sum[49] ^carry[49];
assign Sum[50]= x_sum[50] ^carry[50];
assign Sum[51]= x_sum[51] ^carry[51];
assign Sum[52]= x_sum[52] ^carry[52];
assign Sum[53]= x_sum[53] ^carry[53];
assign Sum[54]= x_sum[54] ^carry[54];
assign Sum[55]= x_sum[55] ^carry[55];
assign Sum[56]= x_sum[56] ^carry[56];
assign Sum[57]= x_sum[57] ^carry[57];
assign Sum[58]= x_sum[58] ^carry[58];
assign Sum[59]= x_sum[59] ^carry[59];
assign Sum[60]= x_sum[60] ^carry[60];
assign Sum[61]= x_sum[61] ^carry[61];
assign Sum[62]= x_sum[62] ^carry[62];
assign Sum[63]= x_sum[63] ^carry[63];
assign Sum[64]= carry[64];


endmodule

module KGP(A,B,kgp);
input [1:0]A,B;
inout [1:0] kgp;
assign kgp[1] = A[1]&A[0] | B[1]&A[0] | A[1]&B[1];
assign kgp[0] = A[1]&A[0] | B[0]&A[0] | A[1]&B[0];
endmodule